library verilog;
use verilog.vl_types.all;
entity EightBitAdder_vlg_vec_tst is
end EightBitAdder_vlg_vec_tst;
