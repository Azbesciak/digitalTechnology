library verilog;
use verilog.vl_types.all;
entity SeqSideEightBitAdder_vlg_vec_tst is
end SeqSideEightBitAdder_vlg_vec_tst;
