library verilog;
use verilog.vl_types.all;
entity FourBitMultiplier_vlg_vec_tst is
end FourBitMultiplier_vlg_vec_tst;
