library verilog;
use verilog.vl_types.all;
entity SeqEightBitAdder_vlg_vec_tst is
end SeqEightBitAdder_vlg_vec_tst;
